module SpecializedMux(I_AM_OWNERS,IRDYS,FRAMES,GLOBAL_IRDY,GLOBAL_FRAME);


input [7:0] I_AM_OWNERS,IRDYS,FRAMES;
output wire GLOBAL_IRDY,GLOBAL_FRAME;

assign {GLOBAL_IRDY,GLOBAL_FRAME} = 
(I_AM_OWNERS[0]) ? {IRDYS[0],FRAMES[0]} :
(I_AM_OWNERS[1]) ? {IRDYS[1],FRAMES[1]} :
(I_AM_OWNERS[2]) ? {IRDYS[2],FRAMES[2]} :
(I_AM_OWNERS[3]) ? {IRDYS[3],FRAMES[3]} :
(I_AM_OWNERS[4]) ? {IRDYS[4],FRAMES[4]} :
(I_AM_OWNERS[5]) ? {IRDYS[5],FRAMES[5]} :
(I_AM_OWNERS[6]) ? {IRDYS[6],FRAMES[6]} :
(I_AM_OWNERS[7]) ? {IRDYS[7],FRAMES[7]} : {1'b1,1'b1};//



endmodule
